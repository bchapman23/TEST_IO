`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:03:00 09/20/2017 
// Design Name: 
// Module Name:    Reveal_Top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////


module Reveal_Top
# (
    parameter NUM_ROWS = 140
)
(
	input  wire [4:0]   okUH,
	output wire [2:0]   okHU,
	inout  wire [31:0]  okUHU,
	inout  wire         okAA,

	input  wire         sys_clk_p,
	input  wire         sys_clk_n,
	
	output wire [7:0]   led,
/*
	inout  wire [31:0]  ddr3_dq,
	output wire [14:0]  ddr3_addr,
	output wire [2 :0]  ddr3_ba,
	output wire [0 :0]  ddr3_ck_p,
	output wire [0 :0]  ddr3_ck_n,
	output wire [0 :0]  ddr3_cke,
	output wire         ddr3_cas_n,
	output wire         ddr3_ras_n,
	output wire         ddr3_we_n,
	output wire [0 :0]  ddr3_odt,
	output wire [3 :0]  ddr3_dm,
	inout  wire [3 :0]  ddr3_dqs_p,
	inout  wire [3 :0]  ddr3_dqs_n,
	output wire         ddr3_reset_n,
*/
	
	/*
	// power spi
	output wire ADC_SYNC1,
	output wire ADC_SYNC2,
	output wire SPI_DI,
	input  wire SPI_DO,
	output wire SPICLK,
	
	// imager spi START HERE
    output wire DIN_T3,
    output wire SPICLK_T3,
    
    // LASER SIGNALS (ignore)
    output wire LE,
    output wire sck,
    output wire mosi,
    output wire ss,
    
    //GALVOs laser and cam (ignore)
    output wire SRI_laser,
    output wire DAC_CLK_laser,
    output wire DAC_LD_n_laser,
    output wire SRI_cam,
    output wire DAC_CLK_cam,
    output wire DAC_LD_n_cam,

    output wire RST_N,
    output wire RS_POT,

    output wire EN_STREAM,              //Enable pattern upload (active high), care
    
    // Clock outputs 
    output wire ADCCLK_IN,          //14.286 MHz clock to ADC
    output wire CLKM,                   //200MHz clock to imager, care
    output wire TX_CLK_IN,  // to sensor, 200MHz serializer clock
    //output wire CLK200MHz,              //200MHz clock to imager for timing of the readout 
    
    output wire PIXGLOB_RES,            //
    // Output signal from readout
    output wire [7:0] ROWADD,           //Row address for readout
    output wire PIXLEFTBUCK_SEL,        //Select the left/right bucket, high for reading left bucket
    output wire PIXRES,
    output wire COL_PRECH,
    output wire ADC_EN,
    output wire DATA_LOAD,
    output wire RST_ADC,
    output wire RST_OUTMUX,
    
    output wire MODDEF,
    
    // Output signal from exposure 
    output wire PIXDRAIN,
    output wire EXP,
    output wire PIXTG,
    output wire DES2, //care
    
    // Mask to sensor
    output wire [10:1] mSTREAM, //care about
    
    output wire FPGA_MOD0,
    output wire FPGA_MOD90,
    
    // i/o for ADC Read 
    input wire TX_CLK_OUT_0,            //clock generated by ADC channel 1-3
    input wire TX_CLK_OUT_1,        //clock generated by ADC channel 4-6
    input wire TX_CLK_OUT_2,            //clock generated by ADC channel 7-9            
    input wire [8:0] DIGOUT,        //care
    
    input  wire    TestIO_3,
    */
    output wire [6:0] TEST_IO,
    
    
	inout wire         IO_SDA,
	inout wire         IO_SCL,
	
	output wire        SPI_DI,
	input wire         SPI_DO,
	output wire        SCLK
	
   );

wire          clk;
wire          rst;

// Clock wizard for base clock
clk_wiz_0 clock_base (
 // Clock in ports
  .clk_in1_p(sys_clk_p),
  .clk_in1_n(sys_clk_n),
  
  // Clock out ports
  .clk_100(clk)
 );

// Front Panel

// Target interface bus:
wire         okClk;
wire [112:0] okHE;
wire [64:0]  okEH;

wire [31:0] select;
wire [31:0] SPIcmd;
wire [31:0] selectButBetter;
reg [6:0] TestIO_reg;



///////

wire CS_POT2;
wire CS_POT1; //THIS IS AN INPUT BECAUSE W16 ISNT WORKING, this provides high impedance
wire COLLOAD_EN;
wire CS_T3;
	
///////////////////////////////////////////

function [7:0] xem7310_led;
input [7:0] a;
integer i;
begin
	for(i=0; i<8; i=i+1) begin: u
		xem7310_led[i] = (a[i]==1'b1) ? (1'b0) : (1'bz);
	end
end
endfunction

assign led = xem7310_led({select[7:0]});
/*
always @*
begin
    if (select == 1) begin
        TestIO_reg[0] = DIN_T3;
        TestIO_reg[1] = SPICLK_T3;
        TestIO_reg[2] = CS_T3;
        TestIO_reg[3] = 0;
        TestIO_reg[4] = 0;
        TestIO_reg[5] = 0;
        TestIO_reg[6] = 0;
    end else if (select == 2) begin
        TestIO_reg[0] = ADCCLK_IN;
        TestIO_reg[1] = CLKM;
        TestIO_reg[2] = TX_CLK_IN;
        TestIO_reg[3] = PIXGLOB_RES;
        TestIO_reg[4] = ROWADD[7];
        TestIO_reg[5] = 0;
        TestIO_reg[6] = 0;
    end else if (select == 3) begin
        TestIO_reg[0] = ROWADD[0];
        TestIO_reg[1] = ROWADD[1];
        TestIO_reg[2] = ROWADD[2];
        TestIO_reg[3] = ROWADD[3];
        TestIO_reg[4] = ROWADD[4];
        TestIO_reg[5] = ROWADD[5];
        TestIO_reg[6] = ROWADD[6];
    end else if (select == 4) begin
        TestIO_reg[0] = PIXLEFTBUCK_SEL;
        TestIO_reg[1] = PIXRES;
        TestIO_reg[2] = COLLOAD_EN;
        TestIO_reg[3] = COL_PRECH;
        TestIO_reg[4] = ADC_EN;
        TestIO_reg[5] = DATA_LOAD;
        TestIO_reg[6] = RST_ADC;
    end else if (select == 5) begin
        TestIO_reg[0] = RST_OUTMUX;
        TestIO_reg[1] = MODDEF;
        TestIO_reg[2] = PIXDRAIN;
        TestIO_reg[3] = EXP;
        TestIO_reg[4] = PIXTG;
        TestIO_reg[5] = DES2;
        TestIO_reg[6] = 0;
    end else if (select == 6) begin
        TestIO_reg[0] = 0;
        TestIO_reg[1] = mSTREAM[1];
        TestIO_reg[2] = mSTREAM[2];
        TestIO_reg[3] = mSTREAM[3];
        TestIO_reg[4] = mSTREAM[4];
        TestIO_reg[5] = mSTREAM[5];
        TestIO_reg[6] = mSTREAM[6];
    end else if (select == 7) begin
        TestIO_reg[0] = mSTREAM[7];
        TestIO_reg[1] = mSTREAM[8];
        TestIO_reg[2] = mSTREAM[9];
        TestIO_reg[3] = mSTREAM[10];
        TestIO_reg[4] = FPGA_MOD0;
        TestIO_reg[5] = FPGA_MOD90;
        TestIO_reg[6] = 0;
    end else if (select == 8) begin
        TestIO_reg[0] = TX_CLK_OUT_0;
        TestIO_reg[1] = TX_CLK_OUT_1;
        TestIO_reg[2] = TX_CLK_OUT_2;
        TestIO_reg[3] = DIGOUT[7];
        TestIO_reg[4] = DIGOUT[8];
        TestIO_reg[5] = TestIO_3;
        TestIO_reg[6] = 0;
    end else if (select == 9) begin
        TestIO_reg[0] = DIGOUT[0];
        TestIO_reg[1] = DIGOUT[1];
        TestIO_reg[2] = DIGOUT[2];
        TestIO_reg[3] = DIGOUT[3];
        TestIO_reg[4] = DIGOUT[4];
        TestIO_reg[5] = DIGOUT[5];
        TestIO_reg[6] = DIGOUT[6];
    end    
end
*/

// Instantiate the okHost and connect endpoints.
wire [65*1-1:0]  okEHx;

okHost okHI(
	.okUH(okUH),
	.okHU(okHU),
	.okUHU(okUHU),
	.okAA(okAA),
	.okClk(okClk),
	.okHE(okHE),
	.okEH(okEH)
	);
                                         
okWireOR # (.N(1)) wireOR (okEH, okEHx);

okWireIn    wi00 (.okHE(okHE),   .ep_addr(8'h00), .ep_dataout(select));  // select


////////////////////////////////////////////////////////
// SPI Test module

// Conditioning to only send instructions when new
reg [31:0] prevData = 32'h0000_0000;
wire newData;
assign newData = (prevData != select);

localparam division = 50;
reg dividedClk = 0;
reg [7:0] subCount = division;
always @ (posedge clk) begin 

    if (subCount == 0) begin 
        dividedClk <= !dividedClk;
        subCount <= division;
        
        
    end else begin
        subCount <= subCount - 1;
        
        // Only update when high following a clock edge
        if ((dividedClk == 1'b1) && (subCount == division)) prevData <= select;
    end
    
end

wire valid;
wire [15:0] CS_STATES;

spi_master_I2Cinterface SPItest(
	.rst(1'b0),
	.clk(clk),
	.wr_clk(dividedClk),
	.wr_en(newData),
	.wr_data(select),
	.busy(i2cBusy),

	.MISO(SPI_DO),	// not enabled
	.MOSI(SPI_DI),
	.SPI_CLK(SCLK),
	.SPI_SS(CS_STATES),
	.valid(valid)
);



///////////////////////////////////////////////////////////
// I2C Code

wire i2cBusy;

i2c_operator # (
    .DIVISION(16'd85) // PCA5555 I/O expanders used can support up to 400 kHz I2C speeds
) i2cSystem (
    .clk(clk),
    .CS(CS_STATES[11:0]),
    .SH_R(6'b0),
    .EN(5'b01100),
    .MUX(1'b0),
    .RS(1'b1),
    .TESTIO(3'b000),

    .reset(1'b0),

    // I2C interface
    .io_sda(IO_SDA),
    .io_scl(IO_SCL),

    .busyI2C(i2cBusy)
);

assign TEST_IO[0] = i2cBusy;
assign TEST_IO[1] = SPI_DO;
assign TEST_IO[2] = SPI_DI;
assign TEST_IO[3] = SCLK;
assign TEST_IO[4] = newData;
assign TEST_IO[5] = valid;
assign TEST_IO[6] = CS_STATES[8];
endmodule
